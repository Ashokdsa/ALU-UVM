`ifndef DWIDTH
  `define DWIDTH 8
  `define CWIDTH 4
  `define LOG2 3
`endif
